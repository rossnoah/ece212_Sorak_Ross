//--------------------------------------------------------------------
// signext.sv - 16-32 bit sign extneder
// David_Harris@hmc.edu 23 October 2005
// Updated to SystemVerilog dmh 12 November 2010
// Refactored into separate files & updated using additional SystemVerilog
// features by John Nestor May 2018
//--------------------------------------------------------------------


module signext(
    input  logic [15:0] a,
    output logic [31:0] y
    );

    assign y = {{16{a[15]}}, a};

endmodule // signext
