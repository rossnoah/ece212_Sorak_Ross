module lab2top (
    ports
);
    
endmodule